library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SinWaveGenerator is
    Port (
        clk : in STD_LOGIC;
        reset : in STD_LOGIC;
        freq : in STD_LOGIC_VECTOR(9 downto 0);
        sync_in : in STD_LOGIC;
        sin_out : out STD_LOGIC_VECTOR(11 downto 0);
        square_out : out STD_LOGIC
    );
end SinWaveGenerator;

architecture Behavioral of SinWaveGenerator is
    signal counter : STD_LOGIC_VECTOR(9 downto 0) := (others => '0');
    signal phase_accumulator : STD_LOGIC_VECTOR(11 downto 0) := (others => '0');  -- Use 12 bits for phase accumulator
    signal rom_address : STD_LOGIC_VECTOR(11 downto 0) := (others => '0');
    signal sine_table : STD_LOGIC_VECTOR(11 downto 0);
    signal sync_edge : STD_LOGIC := '0';

    type ROM is array (0 to 180) of STD_LOGIC_VECTOR(11 downto 0);
    constant sine_rom : ROM := (
        "000000000000",
"000000100011",
"000001000111",
"000001101011",
"000010001110",
"000010110010",
"000011010101",
"000011111001",
"000100011100",
"000101000000",
"000101100011",
"000110000110",
"000110101001",
"000111001100",
"000111101111",
"001000010001",
"001000110100",
"001001010110",
"001001111000",
"001010011010",
"001010111100",
"001011011101",
"001011111110",
"001100011111",
"001101000000",
"001101100001",
"001110000001",
"001110100001",
"001111000001",
"001111100000",
"001111111111",
"010000011110",
"010000111100",
"010001011010",
"010001111000",
"010010010110",
"010010110011",
"010011001111",
"010011101100",
"010100001000",
"010100100011",
"010100111110",
"010101011001",
"010101110100",
"010110001101",
"010110100111",
"010111000000",
"010111011001",
"010111110001",
"011000001000",
"011000100000",
"011000110110",
"011001001101",
"011001100010",
"011001111000",
"011010001100",
"011010100001",
"011010110100",
"011011000111",
"011011011010",
"011011101100",
"011011111110",
"011100001111",
"011100011111",
"011100101111",
"011100111111",
"011101001110",
"011101011100",
"011101101001",
"011101110111",
"011110000011",
"011110001111",
"011110011010",
"011110100101",
"011110101111",
"011110111001",
"011111000010",
"011111001010",
"011111010010",
"011111011001",
"011111011111",
"011111100101",
"011111101011",
"011111101111",
"011111110011",
"011111110111",
"011111111010",
"011111111100",
"011111111101",
"011111111110",
"011111111111",
"011111111110",
"011111111101",
"011111111100",
"011111111010",
"011111110111",
"011111110011",
"011111101111",
"011111101011",
"011111100101",
"011111011111",
"011111011001",
"011111010010",
"011111001010",
"011111000010",
"011110111001",
"011110101111",
"011110100101",
"011110011010",
"011110001111",
"011110000011",
"011101110111",
"011101101001",
"011101011100",
"011101001110",
"011100111111",
"011100101111",
"011100011111",
"011100001111",
"011011111110",
"011011101100",
"011011011010",
"011011000111",
"011010110100",
"011010100001",
"011010001100",
"011001111000",
"011001100010",
"011001001101",
"011000110110",
"011000100000",
"011000001000",
"010111110001",
"010111011001",
"010111000000",
"010110100111",
"010110001101",
"010101110100",
"010101011001",
"010100111110",
"010100100011",
"010100001000",
"010011101100",
"010011001111",
"010010110011",
"010010010110",
"010001111000",
"010001011010",
"010000111100",
"010000011110",
"001111111111",
"001111100000",
"001111000001",
"001110100001",
"001110000001",
"001101100001",
"001101000000",
"001100011111",
"001011111110",
"001011011101",
"001010111100",
"001010011010",
"001001111000",
"001001010110",
"001000110100",
"001000010001",
"000111101111",
"000111001100",
"000110101001",
"000110000110",
"000101100011",
"000101000000",
"000100011100",
"000011111001",
"000011010101",
"000010110010",
"000010001110",
"000001101011",
"000001000111",
"000000100011",
"000000000000"
    );

begin
    process(clk, reset, sync_in)
    begin
        if reset = '1' then
            counter <= (others => '0');
            phase_accumulator <= (others => '0');
            sync_edge <= '0';
        elsif rising_edge(clk) then
            if sync_in = '1' and sync_edge = '0' then
                sync_edge <= '1';
                counter <= (others => '0');
                phase_accumulator <= (others => '0');
            else
                sync_edge <= sync_in;
                counter <= counter + 1;
                if counter = freq then
                    counter <= (others => '0');
                    phase_accumulator <= phase_accumulator + 1;
                    if phase_accumulator = "111111111111" then  -- Adjust the limit for 12 bits
                        phase_accumulator <= (others => '0');
                    end if;
                end if;
            end if;
        end if;
    end process;

    -- ROM lookup
    rom_address <= phase_accumulator;

    -- Create the full sine wave using symmetry
    sine_table <= sine_rom(to_integer(unsigned(rom_address)));
    -- sine_table(11 downto 0) <= sine_table(11 downto 0) & not sine_table(11);  -- Invert the second half

    sin_out <= sine_table;
    square_out <= '1' when phase_accumulator(11) = '1' else '0';

end Behavioral;
